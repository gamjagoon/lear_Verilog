module OR (
input wire A,
input wire B,
output wire C
);

assign C = A | B;

endmodule